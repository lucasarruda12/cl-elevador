library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity floor_checker is
  port (
  );
end floor_checker;

architecture arch of floor_checker is

begin

end arch;